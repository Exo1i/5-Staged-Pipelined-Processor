LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE pkg_opcodes IS
    -- Instruction Opcodes (5-bit)
    CONSTANT OP_NOP : STD_LOGIC_VECTOR(4 DOWNTO 0) := "00000";
    CONSTANT OP_HLT : STD_LOGIC_VECTOR(4 DOWNTO 0) := "00001";
    CONSTANT OP_SETC : STD_LOGIC_VECTOR(4 DOWNTO 0) := "00010";
    CONSTANT OP_NOT : STD_LOGIC_VECTOR(4 DOWNTO 0) := "00011";
    CONSTANT OP_INC : STD_LOGIC_VECTOR(4 DOWNTO 0) := "00100";
    CONSTANT OP_OUT : STD_LOGIC_VECTOR(4 DOWNTO 0) := "00101";
    CONSTANT OP_IN : STD_LOGIC_VECTOR(4 DOWNTO 0) := "00110";
    CONSTANT OP_MOV : STD_LOGIC_VECTOR(4 DOWNTO 0) := "00111";
    CONSTANT OP_SWAP : STD_LOGIC_VECTOR(4 DOWNTO 0) := "01000";
    CONSTANT OP_ADD : STD_LOGIC_VECTOR(4 DOWNTO 0) := "01001";
    CONSTANT OP_SUB : STD_LOGIC_VECTOR(4 DOWNTO 0) := "01010";
    CONSTANT OP_AND : STD_LOGIC_VECTOR(4 DOWNTO 0) := "01011";
    CONSTANT OP_IADD : STD_LOGIC_VECTOR(4 DOWNTO 0) := "01100";
    CONSTANT OP_PUSH : STD_LOGIC_VECTOR(4 DOWNTO 0) := "01101";
    CONSTANT OP_POP : STD_LOGIC_VECTOR(4 DOWNTO 0) := "01110";
    CONSTANT OP_LDM : STD_LOGIC_VECTOR(4 DOWNTO 0) := "01111";
    CONSTANT OP_LDD : STD_LOGIC_VECTOR(4 DOWNTO 0) := "10000";
    CONSTANT OP_STD : STD_LOGIC_VECTOR(4 DOWNTO 0) := "10001";
    CONSTANT OP_JZ : STD_LOGIC_VECTOR(4 DOWNTO 0) := "10010";
    CONSTANT OP_JN : STD_LOGIC_VECTOR(4 DOWNTO 0) := "10011";
    CONSTANT OP_JC : STD_LOGIC_VECTOR(4 DOWNTO 0) := "10100";
    CONSTANT OP_JMP : STD_LOGIC_VECTOR(4 DOWNTO 0) := "10101";
    CONSTANT OP_CALL : STD_LOGIC_VECTOR(4 DOWNTO 0) := "10110";
    CONSTANT OP_RET : STD_LOGIC_VECTOR(4 DOWNTO 0) := "10111";
    CONSTANT OP_INT : STD_LOGIC_VECTOR(4 DOWNTO 0) := "11000";
    CONSTANT OP_RTI : STD_LOGIC_VECTOR(4 DOWNTO 0) := "11001";

    -- Override Operation Types (2-bit)
    CONSTANT OVERRIDE_PUSH_PC : STD_LOGIC_VECTOR(1 DOWNTO 0) := "00";
    CONSTANT OVERRIDE_PUSH_FLAGS : STD_LOGIC_VECTOR(1 DOWNTO 0) := "01";
    CONSTANT OVERRIDE_POP_FLAGS : STD_LOGIC_VECTOR(1 DOWNTO 0) := "10";
    CONSTANT OVERRIDE_POP_PC : STD_LOGIC_VECTOR(1 DOWNTO 0) := "11";

    -- ALU Operations (3-bit)
    CONSTANT ALU_ADD : STD_LOGIC_VECTOR(2 DOWNTO 0) := "000";
    CONSTANT ALU_SUB : STD_LOGIC_VECTOR(2 DOWNTO 0) := "001";
    CONSTANT ALU_AND : STD_LOGIC_VECTOR(2 DOWNTO 0) := "010";
    CONSTANT ALU_NOT : STD_LOGIC_VECTOR(2 DOWNTO 0) := "011";
    CONSTANT ALU_INC : STD_LOGIC_VECTOR(2 DOWNTO 0) := "100";
    CONSTANT ALU_PASS_A : STD_LOGIC_VECTOR(2 DOWNTO 0) := "101";
    CONSTANT ALU_PASS_B : STD_LOGIC_VECTOR(2 DOWNTO 0) := "110";
    CONSTANT ALU_SETC : STD_LOGIC_VECTOR(2 DOWNTO 0) := "111";

    -- OutBSelect Values (2-bit)
    CONSTANT OUTB_REGFILE : STD_LOGIC_VECTOR(1 DOWNTO 0) := "00";
    CONSTANT OUTB_PUSHED_PC : STD_LOGIC_VECTOR(1 DOWNTO 0) := "01";
    CONSTANT OUTB_IMMEDIATE : STD_LOGIC_VECTOR(1 DOWNTO 0) := "10";
    CONSTANT OUTB_INPUT_PORT : STD_LOGIC_VECTOR(1 DOWNTO 0) := "11";

    -- Conditional Types (2-bit)
    CONSTANT COND_ZERO : STD_LOGIC_VECTOR(1 DOWNTO 0) := "00"; -- JZ
    CONSTANT COND_NEGATIVE : STD_LOGIC_VECTOR(1 DOWNTO 0) := "01"; -- JN
    CONSTANT COND_CARRY : STD_LOGIC_VECTOR(1 DOWNTO 0) := "10"; -- JC
    CONSTANT COND_NONE : STD_LOGIC_VECTOR(1 DOWNTO 0) := "11"; -- Unconditional

    -- PassInterrupt Values (2-bit)
    CONSTANT PASS_INT_NORMAL : STD_LOGIC_VECTOR(1 DOWNTO 0) := "00"; -- Normal address from EX/MEM
    CONSTANT PASS_INT_RESET : STD_LOGIC_VECTOR(1 DOWNTO 0) := "01"; -- Reset vector (position 0)
    CONSTANT PASS_INT_SOFTWARE : STD_LOGIC_VECTOR(1 DOWNTO 0) := "10"; -- Software interrupt (from immediate) Immediate + 2
    CONSTANT PASS_INT_HARDWARE : STD_LOGIC_VECTOR(1 DOWNTO 0) := "11"; -- Hardware interrupt (fixed position 1)

    -- Branch Target Select Values (2-bit)
    CONSTANT TARGET_DECODE : STD_LOGIC_VECTOR(1 DOWNTO 0) := "00"; -- Immediate from decode
    CONSTANT TARGET_EXECUTE : STD_LOGIC_VECTOR(1 DOWNTO 0) := "01"; -- Immediate from execute
    CONSTANT TARGET_MEMORY : STD_LOGIC_VECTOR(1 DOWNTO 0) := "10"; -- Interrupt address from memory
    CONSTANT TARGET_RESET : STD_LOGIC_VECTOR(1 DOWNTO 0) := "11"; -- Reset address (0)

    -- Branch Predictor States (2-bit saturating counter)
    CONSTANT STRONGLY_NOT_TAKEN : STD_LOGIC_VECTOR(1 DOWNTO 0) := "00";
    CONSTANT WEAKLY_NOT_TAKEN : STD_LOGIC_VECTOR(1 DOWNTO 0) := "01";
    CONSTANT WEAKLY_TAKEN : STD_LOGIC_VECTOR(1 DOWNTO 0) := "10";
    CONSTANT STRONGLY_TAKEN : STD_LOGIC_VECTOR(1 DOWNTO 0) := "11";

END PACKAGE pkg_opcodes;